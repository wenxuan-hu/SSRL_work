package mc_top_test_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "tb_defs.svh"
    
    `include "dfi_monitor.svh"
    `include "dfi_lpddr4_responder.svh"
    `include "dfi_lpddr4_monitor.svh"
    `include "dfi_lpddr4_agent.svh"

    `include "dla_trans.svh"
    `include "dla_cmd_sequence.svh"
    `include "dla_sequencer.svh"
    `include "dla_driver.svh"
    `include "dla_monitor.svh"
    `include "dla_agent.svh"

    `include "mc_top_checker.svh"
    `include "mc_top_virtual_sequencer.svh"
    `include "mc_top_env.svh"
    `include "mc_top_basic_test.svh"

endpackage
