module mc_core_nointerface_wrapper(

	//system clock/reset
	input clk,
	input rst,

    native_interface native_if_0,
    native_interface native_if_1,
    dfi_lpddr4_interface dfi_lpddr4_if,

    //CSR
    input [1:0] mul_rd_phase_cfg,
    input [1:0] mul_wr_phase_cfg,
    input [1:0] mul_rdcmd_phase_cfg,
    input [1:0] mul_wrcmd_phase_cfg,
    input [7:0] mul_tRRD_cfg,
    input [7:0] mul_tFAW_cfg,
    input [7:0] mul_tCCD_cfg,
    input [7:0] mul_WTR_LATENCY_cfg,
    input [7:0] mul_RTW_LATENCY_cfg,
    input [7:0] mul_READ_TIME_cfg,
    input [7:0] mul_WRITE_TIME_cfg,

    input [11:0] ref_tREFI_cfg,
    input [3:0] ref_POSTPONE_cfg,
    input [7:0] ref_tRP_cfg,
    input [7:0] ref_tRFC_cfg,

    input [7:0] bm_tWTP_cfg,
    input [7:0] bm_tRTP_cfg,
    input [7:0] bm_tRAS_cfg,
    input [7:0] bm_tRC_cfg,
    input [7:0] bm_tRP_cfg,
    input [7:0] bm_tRCD_cfg,
    input [7:0] bm_tCCDMW_cfg,

    input [7:0] crb_READ_LATENCY_cfg,
    input [7:0] crb_WRITE_LATENCY_cfg,
    input [7:0] dfi_rddata_en_latency_cfg,
    input [7:0] dfi_wrdata_en_latency_cfg,

    input [7:0] dfi_wdqs_preamble_cfg
);
mc_core_nointerface u_mc_core_nointerface   (
    .clk	(clk),
	.rst	(rst),

	.mul_rd_phase_cfg	(mul_rd_phase_cfg),
	.mul_wr_phase_cfg	(mul_wr_phase_cfg),
	.mul_rdcmd_phase_cfg	(mul_rdcmd_phase_cfg),
	.mul_wrcmd_phase_cfg	(mul_wrcmd_phase_cfg),
	.mul_tRRD_cfg	(mul_tRRD_cfg),
	.mul_tFAW_cfg	(mul_tFAW_cfg),
	.mul_tCCD_cfg	(mul_tCCD_cfg),
	.mul_WTR_LATENCY_cfg	(mul_WTR_LATENCY_cfg),
	.mul_RTW_LATENCY_cfg	(mul_RTW_LATENCY_cfg),
	.mul_READ_TIME_cfg	(mul_READ_TIME_cfg),
	.mul_WRITE_TIME_cfg (mul_WRITE_TIME_cfg),
	.ref_tREFI_cfg	(ref_tREFI_cfg),
	.ref_POSTPONE_cfg	(ref_POSTPONE_cfg),
	.ref_tRP_cfg	(ref_tRP_cfg),
	.ref_tRFC_cfg	(ref_tRFC_cfg),
	.bm_tWTP_cfg	(bm_tWTP_cfg),
	.bm_tRTP_cfg	(bm_tRTP_cfg),
	.bm_tRAS_cfg	(bm_tRAS_cfg),
	.bm_tRC_cfg		(bm_tRC_cfg),
	.bm_tRP_cfg		(bm_tRP_cfg),
	.bm_tRCD_cfg	(bm_tRCD_cfg),
	.bm_tCCDMW_cfg	(bm_tCCDMW_cfg),
	.crb_READ_LATENCY_cfg	(crb_READ_LATENCY_cfg),
	.crb_WRITE_LATENCY_cfg	(crb_WRITE_LATENCY_cfg),
	.dfi_rddata_en_latency_cfg	(dfi_rddata_en_latency_cfg),
	.dfi_wrdata_en_latency_cfg	(dfi_wrdata_en_latency_cfg),
	.dfi_wdqs_preamble_cfg	(dfi_wdqs_preamble_cfg),
	
	// native interface 0
	.cmd_valid	(native_if_0.native_cmd_valid),
	.cmd_ready	(native_if_0.native_cmd_ready),
	.cmd_first	(native_if_0.native_cmd_first),
	.cmd_last	(native_if_0.native_cmd_last),
	.cmd_payload_we	(native_if_0.native_cmd_payload_we),
	.cmd_payload_mw	(native_if_0.native_cmd_payload_mw),
	.cmd_payload_addr	(native_if_0.native_cmd_payload_addr),
	.wdata_valid	(native_if_0.wdata_valid),
	.wdata_ready	(native_if_0.wdata_ready),
	.wdata_first	(native_if_0.wdata_first),
	.wdata_last		(native_if_0.wdata_last),
	.wdata_payload_data		(native_if_0.wdata_payload_data),
	.wdata_payload_we		(native_if_0.wdata_payload_we),
	.rdata_valid		(native_if_0.rdata_valid),
	.rdata_ready		(native_if_0.rdata_ready),
	.rdata_first		(native_if_0.rdata_first),
	.rdata_last			(native_if_0.rdata_last),
	.rdata_payload_data	(native_if_0.rdata_payload_data),

	// native interface 1
	.cmd_valid_1	(native_if_1.native_cmd_valid),
	.cmd_ready_1	(native_if_1.native_cmd_ready),
	.cmd_first_1	(native_if_1.native_cmd_first),
	.cmd_last_1	(native_if_1.native_cmd_last),
	.cmd_payload_we_1	(native_if_1.native_cmd_payload_we),
	.cmd_payload_mw_1	(native_if_1.native_cmd_payload_mw),
	.cmd_payload_addr_1	(native_if_1.native_cmd_payload_addr),
	.wdata_valid_1	(native_if_1.wdata_valid),
	.wdata_ready_1	(native_if_1.wdata_ready),
	.wdata_first_1	(native_if_1.wdata_first),
	.wdata_last_1		(native_if_1.wdata_last),
	.wdata_payload_data_1		(native_if_1.wdata_payload_data),
	.wdata_payload_we_1		(native_if_1.wdata_payload_we),
	.rdata_valid_1		(native_if_1.rdata_valid),
	.rdata_ready_1		(native_if_1.rdata_ready),
	.rdata_first_1		(native_if_1.rdata_first),
	.rdata_last_1			(native_if_1.rdata_last),
	.rdata_payload_data_1	(native_if_1.rdata_payload_data),
	
	// dfi interface
	.dfi_lpddr4_if_dfi_ca_0	(dfi_lpddr4_if.dfi_phase0_lpddr4_if.ca),
	.dfi_lpddr4_if_dfi_cs_0	(dfi_lpddr4_if.dfi_phase0_lpddr4_if.cs),
	.dfi_lpddr4_if_dfi_cke_0 (dfi_lpddr4_if.dfi_phase0_lpddr4_if.cke),
	.dfi_lpddr4_if_dfi_odt_0 (dfi_lpddr4_if.dfi_phase0_lpddr4_if.odt),
	.dfi_lpddr4_if_dfi_reset_n_0 (dfi_lpddr4_if.dfi_phase0_lpddr4_if.reset_n),
	.dfi_lpddr4_if_dfi_act_n_0	(dfi_lpddr4_if.dfi_phase0_lpddr4_if.act_n),
	.dfi_lpddr4_if_dfi_wrdata_0	(dfi_lpddr4_if.dfi_phase0_lpddr4_if.wrdata),
	.dfi_lpddr4_if_dfi_wrdata_mask_0 (dfi_lpddr4_if.dfi_phase0_lpddr4_if.wrdata_mask),
	.dfi_lpddr4_if_dfi_rdata_0	(dfi_lpddr4_if.dfi_phase0_lpddr4_if.rddata),
	.dfi_lpddr4_if_dfi_rddata_valid_0	(dfi_lpddr4_if.dfi_phase0_lpddr4_if.rddata_valid),
	.dfi_lpddr4_if_dfi_rddata_en_0	(dfi_lpddr4_if.dfi_phase0_lpddr4_if.rddata_en),
	.dfi_lpddr4_if_dfi_wrdata_en_0 (dfi_lpddr4_if.dfi_phase0_lpddr4_if.wrdata_en),

	
	.dfi_lpddr4_if_dfi_ca_1	(dfi_lpddr4_if.dfi_phase1_lpddr4_if.ca),
	.dfi_lpddr4_if_dfi_cs_1 	(dfi_lpddr4_if.dfi_phase1_lpddr4_if.cs),
	.dfi_lpddr4_if_dfi_cke_1 (dfi_lpddr4_if.dfi_phase1_lpddr4_if.cke),
	.dfi_lpddr4_if_dfi_odt_1 (dfi_lpddr4_if.dfi_phase1_lpddr4_if.odt),
	.dfi_lpddr4_if_dfi_reset_n_1 (dfi_lpddr4_if.dfi_phase1_lpddr4_if.reset_n),
	.dfi_lpddr4_if_dfi_act_n_1	(dfi_lpddr4_if.dfi_phase1_lpddr4_if.act_n),
	.dfi_lpddr4_if_dfi_wrdata_1	(dfi_lpddr4_if.dfi_phase1_lpddr4_if.wrdata),
	.dfi_lpddr4_if_dfi_wrdata_mask_1 (dfi_lpddr4_if.dfi_phase1_lpddr4_if.wrdata_mask),
	.dfi_lpddr4_if_dfi_rdata_1	(dfi_lpddr4_if.dfi_phase1_lpddr4_if.rddata),
	.dfi_lpddr4_if_dfi_rddata_valid_1	(dfi_lpddr4_if.dfi_phase1_lpddr4_if.rddata_valid),
	.dfi_lpddr4_if_dfi_rddata_en_1	(dfi_lpddr4_if.dfi_phase1_lpddr4_if.rddata_en),
	.dfi_lpddr4_if_dfi_wrdata_en_1 (dfi_lpddr4_if.dfi_phase1_lpddr4_if.wrdata_en),


	.dfi_lpddr4_if_dfi_ca_2	(dfi_lpddr4_if.dfi_phase2_lpddr4_if.ca),
	.dfi_lpddr4_if_dfi_cs_2 	(dfi_lpddr4_if.dfi_phase2_lpddr4_if.cs),
	.dfi_lpddr4_if_dfi_cke_2 (dfi_lpddr4_if.dfi_phase2_lpddr4_if.cke),
	.dfi_lpddr4_if_dfi_odt_2 (dfi_lpddr4_if.dfi_phase2_lpddr4_if.odt),
	.dfi_lpddr4_if_dfi_reset_n_2 (dfi_lpddr4_if.dfi_phase2_lpddr4_if.reset_n),
	.dfi_lpddr4_if_dfi_act_n_2	(dfi_lpddr4_if.dfi_phase2_lpddr4_if.act_n),
	.dfi_lpddr4_if_dfi_wrdata_2	(dfi_lpddr4_if.dfi_phase2_lpddr4_if.wrdata),
	.dfi_lpddr4_if_dfi_wrdata_mask_2 (dfi_lpddr4_if.dfi_phase2_lpddr4_if.wrdata_mask),
	.dfi_lpddr4_if_dfi_rdata_2	(dfi_lpddr4_if.dfi_phase2_lpddr4_if.rddata),
	.dfi_lpddr4_if_dfi_rddata_valid_2	(dfi_lpddr4_if.dfi_phase2_lpddr4_if.rddata_valid),
	.dfi_lpddr4_if_dfi_rddata_en_2	(dfi_lpddr4_if.dfi_phase2_lpddr4_if.rddata_en),
	.dfi_lpddr4_if_dfi_wrdata_en_2 (dfi_lpddr4_if.dfi_phase2_lpddr4_if.wrdata_en),


	.dfi_lpddr4_if_dfi_ca_3	(dfi_lpddr4_if.dfi_phase3_lpddr4_if.ca),
	.dfi_lpddr4_if_dfi_cs_3 	(dfi_lpddr4_if.dfi_phase3_lpddr4_if.cs),
	.dfi_lpddr4_if_dfi_cke_3 (dfi_lpddr4_if.dfi_phase3_lpddr4_if.cke),
	.dfi_lpddr4_if_dfi_odt_3 (dfi_lpddr4_if.dfi_phase3_lpddr4_if.odt),
	.dfi_lpddr4_if_dfi_reset_n_3 (dfi_lpddr4_if.dfi_phase3_lpddr4_if.reset_n),
	.dfi_lpddr4_if_dfi_act_n_3	(dfi_lpddr4_if.dfi_phase3_lpddr4_if.act_n),
	.dfi_lpddr4_if_dfi_wrdata_3	(dfi_lpddr4_if.dfi_phase3_lpddr4_if.wrdata),
	.dfi_lpddr4_if_dfi_wrdata_mask_3 (dfi_lpddr4_if.dfi_phase3_lpddr4_if.wrdata_mask),
	.dfi_lpddr4_if_dfi_rdata_3	(dfi_lpddr4_if.dfi_phase3_lpddr4_if.rddata),
	.dfi_lpddr4_if_dfi_rddata_valid_3	(dfi_lpddr4_if.dfi_phase3_lpddr4_if.rddata_valid),
	.dfi_lpddr4_if_dfi_rddata_en_3	(dfi_lpddr4_if.dfi_phase3_lpddr4_if.rddata_en),
	.dfi_lpddr4_if_dfi_wrdata_en_3 (dfi_lpddr4_if.dfi_phase3_lpddr4_if.wrdata_en)
	
);

endmodule
