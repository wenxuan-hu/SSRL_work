package ucie_channel_test_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "tb_defs.svh"

    `include "rdi_mb_trans.svh"
    `include "rdi_mb_sequence.svh"
    `include "rdi_mb_sequencer.svh"
    `include "rdi_mb_driver.svh"
    `include "rdi_mb_monitor.svh"
    `include "rdi_mb_agent.svh"

    `include "ucie_channel_checker.svh"
    `include "ucie_channel_virtual_sequencer.svh"
    `include "ucie_channel_env.svh"
    `include "ucie_channel_basic_test.svh"

endpackage