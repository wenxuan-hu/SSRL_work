module  ucie();






endmodule
