package bank_machine_test_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "tb_defs.svh"
    `include "dfi_lpddr4_monitor.svh"

    `include "dfi_trans.svh"
    `include "dfi_cmd_sequence.svh"
    `include "dfi_sequencer.svh"
    `include "dfi_driver.svh"
    `include "dfi_monitor.svh"
    `include "dfi_agent.svh"

    //`include "bm_responder.svh"
    `include "DFIAdapter_checker.svh"
    `include "DFIAdapter_virtual_sequencer.svh"
    `include "DFIAdapter_env.svh"
    `include "DFIAdapter_basic_test.svh"

endpackage