interface top_interface;
// ----------------------------------------------------
//input
    logic             clk  ;
    logic             rst_n  ;
    //TODO   clock and reset signal need to be separated;






      
//clocking drv_cb @(posedge clk);
//default input #10ns output #5ns;
//    output             clk,rst   ;
//    input           rd_ready_o;
//endclocking
//
//clocking mon_cb @(posedge clk);
//default input #10ns output #5ns;
//    input           rd_i;
//
//
//endclocking
      
//modport (input  a, b, output c,d);




endinterface
