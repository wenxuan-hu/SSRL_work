module bankmachine_wrapper(input clk,rst,
    litedram_interface litedram_if,
    cmd_rw_interface cmd_rw_if_0,
    cmd_rw_interface cmd_rw_if_1,
    cmd_rw_interface cmd_rw_if_2,
    cmd_rw_interface cmd_rw_if_3,
    cmd_rw_interface cmd_rw_if_4,
    cmd_rw_interface cmd_rw_if_5,
    cmd_rw_interface cmd_rw_if_6,
    cmd_rw_interface cmd_rw_if_7,
    input [7:0] bm_tRTP_cfg,
	input [7:0] bm_tWTP_cfg,
	input [7:0] bm_tRC_cfg,
	input [7:0] bm_tRAS_cfg,
	input [7:0] bm_tRP_cfg,
	input [7:0] bm_tRCD_cfg,
	input [7:0] bm_tCCDMW_cfg
);
    bankmachine_0 u_bankmachine_0 (
    .req_valid               (litedram_if.litedram_cmd_if_0.interface_bank_valid),
    .req_ready               (litedram_if.litedram_cmd_if_0.interface_bank_ready),
    .req_mw                  (litedram_if.litedram_cmd_if_0.interface_bank_mw),
    .req_we                  (litedram_if.litedram_cmd_if_0.interface_bank_we),
    .req_addr                (litedram_if.litedram_cmd_if_0.interface_bank_addr),
    .req_lock                (litedram_if.litedram_cmd_if_0.interface_bank_lock),
    .req_wdata_ready         (litedram_if.litedram_cmd_if_0.interface_bank_wdata_ready),
    .req_rdata_valid         (litedram_if.litedram_cmd_if_0.interface_bank_rdata_valid),
    .refresh_req             (cmd_rw_if_0.refresh_req),
    .refresh_gnt             (cmd_rw_if_0.refresh_gnt),
    .cmd_valid               (cmd_rw_if_0.cmd_valid),
    .cmd_ready               (cmd_rw_if_0.cmd_ready),
    .cmd_first               (cmd_rw_if_0.cmd_first),
    .cmd_last                (cmd_rw_if_0.cmd_last),
    .cmd_payload_a           (cmd_rw_if_0.cmd_payload_a),
    .cmd_payload_ba          (cmd_rw_if_0.cmd_payload_ba),
    .cmd_payload_cas         (cmd_rw_if_0.cmd_payload_cas),
    .cmd_payload_ras         (cmd_rw_if_0.cmd_payload_ras),
    .cmd_payload_we          (cmd_rw_if_0.cmd_payload_we),
    .cmd_payload_is_cmd      (cmd_rw_if_0.cmd_payload_is_cmd),
    .cmd_payload_is_read     (cmd_rw_if_0.cmd_payload_is_read),
    .cmd_payload_is_write    (cmd_rw_if_0.cmd_payload_is_write),
    .cmd_payload_is_mw       (cmd_rw_if_0.cmd_payload_is_mw),
    .bm_tRTP_cfg             (bm_tRTP_cfg),
    .bm_tWTP_cfg             (bm_tWTP_cfg),
    .bm_tRC_cfg              (bm_tRC_cfg),
    .bm_tRAS_cfg             (bm_tRAS_cfg),
    .bm_tRP_cfg              (bm_tRP_cfg),
    .bm_tRCD_cfg             (bm_tRCD_cfg),
    .bm_tCCDMW_cfg           (bm_tCCDMW_cfg),
    .sys_clk                 (clk),
    .sys_rst                 (rst)
);

    bankmachine_1 u_bankmachine_1 (
    .req_valid               (litedram_if.litedram_cmd_if_1.interface_bank_valid),
    .req_ready               (litedram_if.litedram_cmd_if_1.interface_bank_ready),
    .req_mw                  (litedram_if.litedram_cmd_if_1.interface_bank_mw),
    .req_we                  (litedram_if.litedram_cmd_if_1.interface_bank_we),
    .req_addr                (litedram_if.litedram_cmd_if_1.interface_bank_addr),
    .req_lock                (litedram_if.litedram_cmd_if_1.interface_bank_lock),
    .req_wdata_ready         (litedram_if.litedram_cmd_if_1.interface_bank_wdata_ready),
    .req_rdata_valid         (litedram_if.litedram_cmd_if_1.interface_bank_rdata_valid),
    .refresh_req             (cmd_rw_if_1.refresh_req),
    .refresh_gnt             (cmd_rw_if_1.refresh_gnt),
    .cmd_valid               (cmd_rw_if_1.cmd_valid),
    .cmd_ready               (cmd_rw_if_1.cmd_ready),
    .cmd_first               (cmd_rw_if_1.cmd_first),
    .cmd_last                (cmd_rw_if_1.cmd_last),
    .cmd_payload_a           (cmd_rw_if_1.cmd_payload_a),
    .cmd_payload_ba          (cmd_rw_if_1.cmd_payload_ba),
    .cmd_payload_cas         (cmd_rw_if_1.cmd_payload_cas),
    .cmd_payload_ras         (cmd_rw_if_1.cmd_payload_ras),
    .cmd_payload_we          (cmd_rw_if_1.cmd_payload_we),
    .cmd_payload_is_cmd      (cmd_rw_if_1.cmd_payload_is_cmd),
    .cmd_payload_is_read     (cmd_rw_if_1.cmd_payload_is_read),
    .cmd_payload_is_write    (cmd_rw_if_1.cmd_payload_is_write),
    .cmd_payload_is_mw       (cmd_rw_if_1.cmd_payload_is_mw),
    .bm_tRTP_cfg             (bm_tRTP_cfg),
    .bm_tWTP_cfg             (bm_tWTP_cfg),
    .bm_tRC_cfg              (bm_tRC_cfg),
    .bm_tRAS_cfg             (bm_tRAS_cfg),
    .bm_tRP_cfg              (bm_tRP_cfg),
    .bm_tRCD_cfg             (bm_tRCD_cfg),
    .bm_tCCDMW_cfg           (bm_tCCDMW_cfg),
    .sys_clk                 (clk),
    .sys_rst                 (rst)
);

    bankmachine_2 u_bankmachine_2 (
    .req_valid               (litedram_if.litedram_cmd_if_2.interface_bank_valid),
    .req_ready               (litedram_if.litedram_cmd_if_2.interface_bank_ready),
    .req_mw                  (litedram_if.litedram_cmd_if_2.interface_bank_mw),
    .req_we                  (litedram_if.litedram_cmd_if_2.interface_bank_we),
    .req_addr                (litedram_if.litedram_cmd_if_2.interface_bank_addr),
    .req_lock                (litedram_if.litedram_cmd_if_2.interface_bank_lock),
    .req_wdata_ready         (litedram_if.litedram_cmd_if_2.interface_bank_wdata_ready),
    .req_rdata_valid         (litedram_if.litedram_cmd_if_2.interface_bank_rdata_valid),
    .refresh_req             (cmd_rw_if_2.refresh_req),
    .refresh_gnt             (cmd_rw_if_2.refresh_gnt),
    .cmd_valid               (cmd_rw_if_2.cmd_valid),
    .cmd_ready               (cmd_rw_if_2.cmd_ready),
    .cmd_first               (cmd_rw_if_2.cmd_first),
    .cmd_last                (cmd_rw_if_2.cmd_last),
    .cmd_payload_a           (cmd_rw_if_2.cmd_payload_a),
    .cmd_payload_ba          (cmd_rw_if_2.cmd_payload_ba),
    .cmd_payload_cas         (cmd_rw_if_2.cmd_payload_cas),
    .cmd_payload_ras         (cmd_rw_if_2.cmd_payload_ras),
    .cmd_payload_we          (cmd_rw_if_2.cmd_payload_we),
    .cmd_payload_is_cmd      (cmd_rw_if_2.cmd_payload_is_cmd),
    .cmd_payload_is_read     (cmd_rw_if_2.cmd_payload_is_read),
    .cmd_payload_is_write    (cmd_rw_if_2.cmd_payload_is_write),
    .cmd_payload_is_mw       (cmd_rw_if_2.cmd_payload_is_mw),
    .bm_tRTP_cfg             (bm_tRTP_cfg),
    .bm_tWTP_cfg             (bm_tWTP_cfg),
    .bm_tRC_cfg              (bm_tRC_cfg),
    .bm_tRAS_cfg             (bm_tRAS_cfg),
    .bm_tRP_cfg              (bm_tRP_cfg),
    .bm_tRCD_cfg             (bm_tRCD_cfg),
    .bm_tCCDMW_cfg           (bm_tCCDMW_cfg),
    .sys_clk                 (clk),
    .sys_rst                 (rst)
);

    bankmachine_3 u_bankmachine_3 (
    .req_valid               (litedram_if.litedram_cmd_if_3.interface_bank_valid),
    .req_ready               (litedram_if.litedram_cmd_if_3.interface_bank_ready),
    .req_mw                  (litedram_if.litedram_cmd_if_3.interface_bank_mw),
    .req_we                  (litedram_if.litedram_cmd_if_3.interface_bank_we),
    .req_addr                (litedram_if.litedram_cmd_if_3.interface_bank_addr),
    .req_lock                (litedram_if.litedram_cmd_if_3.interface_bank_lock),
    .req_wdata_ready         (litedram_if.litedram_cmd_if_3.interface_bank_wdata_ready),
    .req_rdata_valid         (litedram_if.litedram_cmd_if_3.interface_bank_rdata_valid),
    .refresh_req             (cmd_rw_if_3.refresh_req),
    .refresh_gnt             (cmd_rw_if_3.refresh_gnt),
    .cmd_valid               (cmd_rw_if_3.cmd_valid),
    .cmd_ready               (cmd_rw_if_3.cmd_ready),
    .cmd_first               (cmd_rw_if_3.cmd_first),
    .cmd_last                (cmd_rw_if_3.cmd_last),
    .cmd_payload_a           (cmd_rw_if_3.cmd_payload_a),
    .cmd_payload_ba          (cmd_rw_if_3.cmd_payload_ba),
    .cmd_payload_cas         (cmd_rw_if_3.cmd_payload_cas),
    .cmd_payload_ras         (cmd_rw_if_3.cmd_payload_ras),
    .cmd_payload_we          (cmd_rw_if_3.cmd_payload_we),
    .cmd_payload_is_cmd      (cmd_rw_if_3.cmd_payload_is_cmd),
    .cmd_payload_is_read     (cmd_rw_if_3.cmd_payload_is_read),
    .cmd_payload_is_write    (cmd_rw_if_3.cmd_payload_is_write),
    .cmd_payload_is_mw       (cmd_rw_if_3.cmd_payload_is_mw),
    .bm_tRTP_cfg             (bm_tRTP_cfg),
    .bm_tWTP_cfg             (bm_tWTP_cfg),
    .bm_tRC_cfg              (bm_tRC_cfg),
    .bm_tRAS_cfg             (bm_tRAS_cfg),
    .bm_tRP_cfg              (bm_tRP_cfg),
    .bm_tRCD_cfg             (bm_tRCD_cfg),
    .bm_tCCDMW_cfg           (bm_tCCDMW_cfg),
    .sys_clk                 (clk),
    .sys_rst                 (rst)
);

    bankmachine_4 u_bankmachine_4 (
    .req_valid               (litedram_if.litedram_cmd_if_4.interface_bank_valid),
    .req_ready               (litedram_if.litedram_cmd_if_4.interface_bank_ready),
    .req_mw                  (litedram_if.litedram_cmd_if_4.interface_bank_mw),
    .req_we                  (litedram_if.litedram_cmd_if_4.interface_bank_we),
    .req_addr                (litedram_if.litedram_cmd_if_4.interface_bank_addr),
    .req_lock                (litedram_if.litedram_cmd_if_4.interface_bank_lock),
    .req_wdata_ready         (litedram_if.litedram_cmd_if_4.interface_bank_wdata_ready),
    .req_rdata_valid         (litedram_if.litedram_cmd_if_4.interface_bank_rdata_valid),
    .refresh_req             (cmd_rw_if_4.refresh_req),
    .refresh_gnt             (cmd_rw_if_4.refresh_gnt),
    .cmd_valid               (cmd_rw_if_4.cmd_valid),
    .cmd_ready               (cmd_rw_if_4.cmd_ready),
    .cmd_first               (cmd_rw_if_4.cmd_first),
    .cmd_last                (cmd_rw_if_4.cmd_last),
    .cmd_payload_a           (cmd_rw_if_4.cmd_payload_a),
    .cmd_payload_ba          (cmd_rw_if_4.cmd_payload_ba),
    .cmd_payload_cas         (cmd_rw_if_4.cmd_payload_cas),
    .cmd_payload_ras         (cmd_rw_if_4.cmd_payload_ras),
    .cmd_payload_we          (cmd_rw_if_4.cmd_payload_we),
    .cmd_payload_is_cmd      (cmd_rw_if_4.cmd_payload_is_cmd),
    .cmd_payload_is_read     (cmd_rw_if_4.cmd_payload_is_read),
    .cmd_payload_is_write    (cmd_rw_if_4.cmd_payload_is_write),
    .cmd_payload_is_mw       (cmd_rw_if_4.cmd_payload_is_mw),
    .bm_tRTP_cfg             (bm_tRTP_cfg),
    .bm_tWTP_cfg             (bm_tWTP_cfg),
    .bm_tRC_cfg              (bm_tRC_cfg),
    .bm_tRAS_cfg             (bm_tRAS_cfg),
    .bm_tRP_cfg              (bm_tRP_cfg),
    .bm_tRCD_cfg             (bm_tRCD_cfg),
    .bm_tCCDMW_cfg           (bm_tCCDMW_cfg),
    .sys_clk                 (clk),
    .sys_rst                 (rst)
);

    bankmachine_5 u_bankmachine_5 (
    .req_valid               (litedram_if.litedram_cmd_if_5.interface_bank_valid),
    .req_ready               (litedram_if.litedram_cmd_if_5.interface_bank_ready),
    .req_mw                  (litedram_if.litedram_cmd_if_5.interface_bank_mw),
    .req_we                  (litedram_if.litedram_cmd_if_5.interface_bank_we),
    .req_addr                (litedram_if.litedram_cmd_if_5.interface_bank_addr),
    .req_lock                (litedram_if.litedram_cmd_if_5.interface_bank_lock),
    .req_wdata_ready         (litedram_if.litedram_cmd_if_5.interface_bank_wdata_ready),
    .req_rdata_valid         (litedram_if.litedram_cmd_if_5.interface_bank_rdata_valid),
    .refresh_req             (cmd_rw_if_5.refresh_req),
    .refresh_gnt             (cmd_rw_if_5.refresh_gnt),
    .cmd_valid               (cmd_rw_if_5.cmd_valid),
    .cmd_ready               (cmd_rw_if_5.cmd_ready),
    .cmd_first               (cmd_rw_if_5.cmd_first),
    .cmd_last                (cmd_rw_if_5.cmd_last),
    .cmd_payload_a           (cmd_rw_if_5.cmd_payload_a),
    .cmd_payload_ba          (cmd_rw_if_5.cmd_payload_ba),
    .cmd_payload_cas         (cmd_rw_if_5.cmd_payload_cas),
    .cmd_payload_ras         (cmd_rw_if_5.cmd_payload_ras),
    .cmd_payload_we          (cmd_rw_if_5.cmd_payload_we),
    .cmd_payload_is_cmd      (cmd_rw_if_5.cmd_payload_is_cmd),
    .cmd_payload_is_read     (cmd_rw_if_5.cmd_payload_is_read),
    .cmd_payload_is_write    (cmd_rw_if_5.cmd_payload_is_write),
    .cmd_payload_is_mw       (cmd_rw_if_5.cmd_payload_is_mw),
    .bm_tRTP_cfg             (bm_tRTP_cfg),
    .bm_tWTP_cfg             (bm_tWTP_cfg),
    .bm_tRC_cfg              (bm_tRC_cfg),
    .bm_tRAS_cfg             (bm_tRAS_cfg),
    .bm_tRP_cfg              (bm_tRP_cfg),
    .bm_tRCD_cfg             (bm_tRCD_cfg),
    .bm_tCCDMW_cfg           (bm_tCCDMW_cfg),
    .sys_clk                 (clk),
    .sys_rst                 (rst)
);

    bankmachine_6 u_bankmachine_6 (
    .req_valid               (litedram_if.litedram_cmd_if_6.interface_bank_valid),
    .req_ready               (litedram_if.litedram_cmd_if_6.interface_bank_ready),
    .req_mw                  (litedram_if.litedram_cmd_if_6.interface_bank_mw),
    .req_we                  (litedram_if.litedram_cmd_if_6.interface_bank_we),
    .req_addr                (litedram_if.litedram_cmd_if_6.interface_bank_addr),
    .req_lock                (litedram_if.litedram_cmd_if_6.interface_bank_lock),
    .req_wdata_ready         (litedram_if.litedram_cmd_if_6.interface_bank_wdata_ready),
    .req_rdata_valid         (litedram_if.litedram_cmd_if_6.interface_bank_rdata_valid),
    .refresh_req             (cmd_rw_if_6.refresh_req),
    .refresh_gnt             (cmd_rw_if_6.refresh_gnt),
    .cmd_valid               (cmd_rw_if_6.cmd_valid),
    .cmd_ready               (cmd_rw_if_6.cmd_ready),
    .cmd_first               (cmd_rw_if_6.cmd_first),
    .cmd_last                (cmd_rw_if_6.cmd_last),
    .cmd_payload_a           (cmd_rw_if_6.cmd_payload_a),
    .cmd_payload_ba          (cmd_rw_if_6.cmd_payload_ba),
    .cmd_payload_cas         (cmd_rw_if_6.cmd_payload_cas),
    .cmd_payload_ras         (cmd_rw_if_6.cmd_payload_ras),
    .cmd_payload_we          (cmd_rw_if_6.cmd_payload_we),
    .cmd_payload_is_cmd      (cmd_rw_if_6.cmd_payload_is_cmd),
    .cmd_payload_is_read     (cmd_rw_if_6.cmd_payload_is_read),
    .cmd_payload_is_write    (cmd_rw_if_6.cmd_payload_is_write),
    .cmd_payload_is_mw       (cmd_rw_if_6.cmd_payload_is_mw),
    .bm_tRTP_cfg             (bm_tRTP_cfg),
    .bm_tWTP_cfg             (bm_tWTP_cfg),
    .bm_tRC_cfg              (bm_tRC_cfg),
    .bm_tRAS_cfg             (bm_tRAS_cfg),
    .bm_tRP_cfg              (bm_tRP_cfg),
    .bm_tRCD_cfg             (bm_tRCD_cfg),
    .bm_tCCDMW_cfg           (bm_tCCDMW_cfg),
    .sys_clk                 (clk),
    .sys_rst                 (rst)
);

    bankmachine_7 u_bankmachine_7 (
    .req_valid               (litedram_if.litedram_cmd_if_7.interface_bank_valid),
    .req_ready               (litedram_if.litedram_cmd_if_7.interface_bank_ready),
    .req_mw                  (litedram_if.litedram_cmd_if_7.interface_bank_mw),
    .req_we                  (litedram_if.litedram_cmd_if_7.interface_bank_we),
    .req_addr                (litedram_if.litedram_cmd_if_7.interface_bank_addr),
    .req_lock                (litedram_if.litedram_cmd_if_7.interface_bank_lock),
    .req_wdata_ready         (litedram_if.litedram_cmd_if_7.interface_bank_wdata_ready),
    .req_rdata_valid         (litedram_if.litedram_cmd_if_7.interface_bank_rdata_valid),
    .refresh_req             (cmd_rw_if_7.refresh_req),
    .refresh_gnt             (cmd_rw_if_7.refresh_gnt),
    .cmd_valid               (cmd_rw_if_7.cmd_valid),
    .cmd_ready               (cmd_rw_if_7.cmd_ready),
    .cmd_first               (cmd_rw_if_7.cmd_first),
    .cmd_last                (cmd_rw_if_7.cmd_last),
    .cmd_payload_a           (cmd_rw_if_7.cmd_payload_a),
    .cmd_payload_ba          (cmd_rw_if_7.cmd_payload_ba),
    .cmd_payload_cas         (cmd_rw_if_7.cmd_payload_cas),
    .cmd_payload_ras         (cmd_rw_if_7.cmd_payload_ras),
    .cmd_payload_we          (cmd_rw_if_7.cmd_payload_we),
    .cmd_payload_is_cmd      (cmd_rw_if_7.cmd_payload_is_cmd),
    .cmd_payload_is_read     (cmd_rw_if_7.cmd_payload_is_read),
    .cmd_payload_is_write    (cmd_rw_if_7.cmd_payload_is_write),
    .cmd_payload_is_mw       (cmd_rw_if_7.cmd_payload_is_mw),
    .bm_tRTP_cfg             (bm_tRTP_cfg),
    .bm_tWTP_cfg             (bm_tWTP_cfg),
    .bm_tRC_cfg              (bm_tRC_cfg),
    .bm_tRAS_cfg             (bm_tRAS_cfg),
    .bm_tRP_cfg              (bm_tRP_cfg),
    .bm_tRCD_cfg             (bm_tRCD_cfg),
    .bm_tCCDMW_cfg           (bm_tCCDMW_cfg),
    .sys_clk                 (clk),
    .sys_rst                 (rst)
);

endmodule