package multiplexer_test_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "tb_defs.svh"

    `include "bm_trans.svh"
    `include "bm_cmd_sequence.svh"
    `include "bm_sequencer.svh"
    `include "bm_driver.svh"
    `include "bm_monitor.svh"
    `include "bm_agent.svh"

    `include "refresher_monitor.svh"

    `include "dfi_monitor.svh"

    `include "dfi_checker.svh"

    `include "multiplexer_virtual_sequencer.svh"
    `include "multiplexer_env.svh"

    `include "multiplexer_basic_test.svh"

endpackage