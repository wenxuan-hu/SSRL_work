/*********************************************************************************
Copyright (c) 2021 Wavious LLC

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.

*********************************************************************************/

`ifdef SYNTHESIS
`else 
// AMS netlist generated by the AMS Unified netlister
// IC subversion:  IC6.1.8-64b.500.14 
// Xcelium version: 20.09-s003
// Copyright(C) 2005-2009, Cadence Design Systems, Inc
// User: shadzibabic Pid: 13323
// Design library name: wphy_gf12lp_ips_sim_lib
// Design cell name: wphy_sa_4g_2ph_pdly_no_esd_tb
// Design view name: config_vlog
// Solver: Spectre



// HDL file - wphy_gf12lp_ips_lib, wphy_sa_4g_2ph_pdly_no_esd_wphy_nmos_switch, systemVerilog.

// Library - wphy_gf12lp_ips_lib, Cell - wphy_sa_4g_2ph_pdly_no_esd,
//View - schematic
// LAST TIME SAVED: Sep 18 06:58:13 2020
// NETLIST TIME: Nov 22 23:24:06 2020
`timescale 1ps / 1ps 




 

`endif //SYNTHESIS 
module wphy_sa_4g_2ph_pdly_no_esd (d_data_c, d_data_t, d_datab_c, 
    d_datab_t,   d_cal_c, d_cal_dir_c, d_cal_dir_t, d_cal_t, 
    d_clk_c, d_clk_t, d_dly_ctrl_c, d_dly_ctrl_t, d_dly_gear_c, 
    d_dly_gear_t, d_sa_ena, d_sacal_ena, rxin, vref
`ifdef WLOGIC_NO_PG 
`else  
 ,vdda  
 ,vss 
`endif //WLOGIC_NO_PG 
);

`ifdef WLOGIC_NO_PG
wire vdda;
assign vdda=1'b1;
wire vss;
assign vss=1'b0;
`else
inout vdda;
inout vss;
`endif


output  d_data_c, d_data_t, d_datab_c, d_datab_t;



input  d_cal_dir_c, d_cal_dir_t, d_clk_c, d_clk_t, d_sa_ena, 
    d_sacal_ena, rxin, vref;

input [1:0]  d_dly_gear_c;
input [5:0]  d_dly_ctrl_c;
input [1:0]  d_dly_gear_t;
input [3:0]  d_cal_t;
input [3:0]  d_cal_c;
input [5:0]  d_dly_ctrl_t;

`ifdef SYNTHESIS
`else 

integer in_sw;

wphy_sa_4g_2ph_pdly_no_esd_wphy_nmos_switch Iswitch ( .ena(d_sacal_ena), .out(in_sw), .vss(vss), 
    .inp(rxin), .inn(vref));

wphy_sa_4g_2ph_pdly_no_esd_wphy_sa_4g_pdly SNSAMP_T ( .cal(d_cal_t), .vdda(vdda), 
    .dly_gear(d_dly_gear_t), .inn(vref), .inp(in_sw), .ena(d_sa_ena), 
    .qb(d_datab_t), .cal_dir(d_cal_dir_t), .q(d_data_t), .vss(vss), 
    .dly_ctrl(d_dly_ctrl_t), .clk(d_clk_t));

wphy_sa_4g_2ph_pdly_no_esd_wphy_sa_4g_pdly SNSAMP_C ( .cal(d_cal_c), .vdda(vdda), 
    .dly_gear(d_dly_gear_c), .inn(vref), .inp(in_sw), .ena(d_sa_ena), 
    .qb(d_datab_c), .cal_dir(d_cal_dir_c), .q(d_data_c), .vss(vss), 
    .dly_ctrl(d_dly_ctrl_c), .clk(d_clk_c));

`endif //SYNTHESIS 
endmodule
`ifdef SYNTHESIS
`else
// Library - wphy_gf12lp_ips_sim_lib, Cell -
//wphy_sa_4g_2ph_pdly_no_esd_tb, View - schematic
// LAST TIME SAVED: Oct 28 23:48:13 2020
// NETLIST TIME: Nov 22 23:24:06 2020
`timescale 1ps / 1ps 




 




 // END AMS-UNL Netlist

//systemVerilog HDL for "wphy_ips_lib", "wphy_sa_4g_2ph_pdly_no_esd_wphy_sa_4g_pdly" "systemVerilog"


`timescale 1ps/1fs

module wphy_sa_4g_2ph_pdly_no_esd_wphy_sa_4g_pdly ( q, qb, vdda, vss, cal, cal_dir, clk, dly_ctrl, dly_gear,
ena, inn, inp );

  input  [3:0] cal;
  input cal_dir;
  output q;
  inout vdda;
  input ena;
  input  [1:0] dly_gear;   //TODO: add freq check and enable impact
  input clk;
`ifdef WPIN_EN
  input var integer inp;
  input var integer inn;
`else
  input var integer inp;
  input  inn;
`endif
  input  [5:0] dly_ctrl;
  inout vss;
  output qb;


`ifdef WPIN_EN
`elsif WPIN_UART_EN
Wpin_uart_rx Winn(inn);
`endif

wire power_ok;
reg in;
reg out_pre;
real SA_OFFSET =0.0;
real cal_v = 0.0;
real delay_step = 2.5;
real delay_total = 0.0;
reg clk_b_int;
wire clk_int;

assign power_ok = (vdda & ~vss);
initial begin
    if ($value$plusargs("SnsAmp_OFFSET=%f", SA_OFFSET)) begin
        //$display("SnsAmp_OFFSET %f.", SA_OFFSET);
    end

    clk_b_int = ~clk;
    out_pre    <= 1'b0;

   if(ena) begin
    case(dly_gear)
      0: delay_total = 40+6*dly_ctrl;
      1: delay_total = 24+3*dly_ctrl;
      2: delay_total = 18+2*dly_ctrl;
      3: delay_total = 15+1*dly_ctrl;
      default: delay_total = 0.0;
    endcase

      clk_b_int <= #(delay_total) ~clk;
   end
   else
      clk_b_int = 1'b1;

end

always @(clk,dly_ctrl,ena,dly_gear) begin
   if(ena) begin
    case(dly_gear)
      0: delay_total = 40+6*dly_ctrl;
      1: delay_total = 24+3*dly_ctrl;
      2: delay_total = 18+2*dly_ctrl;
      3: delay_total = 15+1*dly_ctrl;
      default: delay_total = 0.0;
    endcase

      clk_b_int <= #(delay_total) ~clk;
   end
   else
      clk_b_int = 1'b1;

end

assign clk_int = ~clk_b_int;

always @(*) begin
  cal_v = 0.0004*(cal)*((-1.0)**cal_dir);
end

real temp;
real temp_2;
real temp_3;

always @(negedge clk_b_int,negedge ena) begin
   if(ena) begin
`ifdef WPIN_EN
      in = (real'(inp)/1000 -real'(inn)/1000 - SA_OFFSET + cal_v)>0;
      if (inp===1'bx | inn===1'bX | inn===1'bZ | inp===1'bZ)
         out_pre <= 1'bx;
      else
         out_pre  <= (real'(inp)/1000 - real'(inn)/1000==SA_OFFSET - cal_v) ? $random : in;
`elsif WPIN_UART_EN
      in = (real'(inp)/1000 -real'(Winn.value)/1000 - SA_OFFSET + cal_v)>0;
      if (inp===1'bx | inn===1'bX | inn===1'bZ | inp===1'bZ)
         out_pre <= 1'bx;
      else
         out_pre  <= (real'(inp)/1000 - real'(Winn.value)/1000==SA_OFFSET - cal_v) ? $random : in;
`else
      //in = (real'(inp)/1000 -real'(inn*500)/1000 - SA_OFFSET + cal_v)>0;
      /*
      temp_2=inp;
      temp_3=inn*500;
      temp=(real'(Iswitch.out)/1000 -real'(inn*500)/1000 - SA_OFFSET + cal_v);
      */
      in = (real'(Iswitch.out)/1000 -real'(inn*500)/1000 - SA_OFFSET + cal_v)>0;
      if (inp===1'bx | inn===1'bX | inn===1'bZ | inp===1'bZ)
         out_pre <= 1'bx;
      else
         //out_pre  <= (real'(inp)/1000 - real'(inn*500)/1000==SA_OFFSET - cal_v) ? $random : in;
         out_pre  <= (real'(Iswitch.out)/1000 - real'(inn*500)/1000==SA_OFFSET - cal_v) ? $random : in;
`endif
   end
   else begin
      out_pre     <= 1'b0;
   end
end


`ifdef SA_BEHAV
assign q = power_ok ? in :1'bx;
`else
assign q = power_ok ? out_pre :1'bx;
`endif
assign qb = power_ok ? ~out_pre :1'bx;


endmodule
//systemVerilog HDL for "wphy_gf12lp_ips_sim_lib", "wphy_real_channel_model"
//"systemVerilog"

`timescale 1ps/1fs
module wphy_sa_4g_2ph_pdly_no_esd_wphy_real_channel_model #(
  parameter     NUM_OF_COEFFS   = 200,
  parameter     TIMESTEP_PS     = 10,
  parameter     COEFF_FILE      = "channel_coeffs_10ps.txt",
  parameter     DELAY           = 0,
  parameter     AMP_RATIO       = 1
)(  rx_in, rxp_out);
 
input   rx_in;

`ifdef WCHANNEL_EN
output var real rxp_out;

var real rxp_out_tmp;
real rx_in_r ;
integer data_file;      //file handler
integer scan_file;      //file handler
integer i;
integer j;
var real tmp_rxp_out;
//parameter real DRV_SUPPLY = 0.4; // but you should use  0.4;
parameter real DRV_SUPPLY = 1.0; // but you should use  0.4;
real chan_coeffs[200];

real coeffs_array[NUM_OF_COEFFS];
real sample_delays[NUM_OF_COEFFS];

real summed_value;

integer skew=0;
integer max_c2c_jit=0;
integer max_accum_jit=0;
integer ration_min=100;
integer ration_max=100;
real    amp_ratio;
wire    rx_in_jitter;

initial begin
  if(rx_in) begin
    rxp_out=1000;
    rxp_out_tmp=1000;
  end
  else begin
    rxp_out=0;
    rxp_out_tmp=0;
  end
end

initial begin
    if ($value$plusargs("RCVR_SKEW=%d", skew)) begin
    end
    if ($value$plusargs("RCVR_MAX_C2C_JIT=%d", max_c2c_jit)) begin
    end
    if ($value$plusargs("RCVR_MAX_ACCUM_JIT=%d", max_accum_jit)) begin
    end
    if ($value$plusargs("RCVR_AMP_RATIO_MIN=%d", ration_min)) begin
    end
    if ($value$plusargs("RCVR_AMP_RATIO_MAX=%d", ration_max)) begin
    end

    amp_ratio=($urandom_range(ration_min,ration_max))/100.0;
end


ddr_jitter_buf u_jitter_buf (
   .i_clk(rx_in),
   .i_skew(skew),
   .i_max_c2c_jit(max_c2c_jit),
   .i_max_accum_jit(max_accum_jit),
   .o_clk(rx_in_jitter)
);

always @(posedge rx_in_jitter) begin
    rxp_out_tmp = 0.0;
  for(j=0;j<5;j=j+1) begin
    #6ps;
    rxp_out_tmp = (200+rxp_out_tmp);
  end
end
always @(negedge rx_in_jitter) begin
    rxp_out_tmp = 1000.0;
  for(j=0;j<5;j=j+1) begin
    #6ps;
    rxp_out_tmp = (rxp_out_tmp-200);
  end
end

always @(rxp_out_tmp) rxp_out=rxp_out_tmp*amp_ratio;

//always @(*) begin 
//   if (rx_in === 1'bz) rx_in_r = 1.234e6;
//   else rx_in_r = (rx_in) ? 1.0 : 0.0;
//end
//
////Coeff math
////Delays go 0 -> NUM_OF_COEFFS
//always #(TIMESTEP_PS) begin
//  summed_value = 0;
//  
//  //Delays
//  for(i=NUM_OF_COEFFS-1; i >=0; i--) begin
//    if(i == 0) begin                //First one is the input 
//      sample_delays[i] = rx_in_r;
//    end else begin                  //remainder are last one
//      sample_delays[i] = sample_delays[i-1];      
//    end
//  end
//  
//  
//  for(i=0; i<NUM_OF_COEFFS; i++) begin
//    //summed_value += coeffs_array[i] * sample_delays[i]; 
//    //summed_value += (chan_coeffs[i]/0.36) * sample_delays[i]; 
//    summed_value += (chan_coeffs[i]/0.15) * sample_delays[i]; 
//  end 
//
//end
//
////assign rxp_out = (rx_in!==1'bz) ? summed_value * DRV_SUPPLY : 1.234e6;
//assign rxp_out_tmp = (rx_in!==1'bz) ? summed_value * DRV_SUPPLY : 1.234e6;
//
//always @(rxp_out_tmp) begin
//       rxp_out <= #(DELAY) rxp_out_tmp*AMP_RATIO;
//end
//
////initial begin  
////  foreach (coeffs_array[i]) begin
////    coeffs_array[i] = chan_coeffs[i]/0.8;
////  end
////end
//
//
////assign chan_coeffs[0] = 0;
////assign chan_coeffs[1] = 0;
////assign chan_coeffs[2] = 0;
////assign chan_coeffs[3] = 0;
////assign chan_coeffs[4] = 0.01;
////assign chan_coeffs[5] = 0.02;
////assign chan_coeffs[6] = 0.03;
////assign chan_coeffs[7] = 0.04;
////assign chan_coeffs[8] = 0.05;
////assign chan_coeffs[9] = 0.05;
////assign chan_coeffs[10] = 0.04;
////assign chan_coeffs[11] = 0.03;
////assign chan_coeffs[12] = 0.02;
////assign chan_coeffs[13] = 0.01;
////assign chan_coeffs[14] = 0.01;
////assign chan_coeffs[15] = 0.01;
////assign chan_coeffs[16] = 0.01;
////assign chan_coeffs[17] = 0.01;
////assign chan_coeffs[18] = 0.01;
////assign chan_coeffs[19] = 0.01;
//
//assign chan_coeffs[0] = 0;
//assign chan_coeffs[1] = 0.02;
//assign chan_coeffs[2] = 0.04;
//assign chan_coeffs[3] = 0.05;
//assign chan_coeffs[4] = 0.03;
//assign chan_coeffs[5] = 0.01;
////assign chan_coeffs[6] = 0.01;
////assign chan_coeffs[7] = 0.01;
////assign chan_coeffs[8] = 0.03;
////assign chan_coeffs[9] = 0.02;
////assign chan_coeffs[10] = 0.04*3;
////assign chan_coeffs[11] = 0.03*3;
////assign chan_coeffs[12] = 0.02*3;
////assign chan_coeffs[13] = 0.01*3;
////assign chan_coeffs[14] = 0.01*3;
////assign chan_coeffs[15] = 0.01*3;
////assign chan_coeffs[16] = 0.01*3;
////assign chan_coeffs[17] = 0.01*3;
////assign chan_coeffs[18] = 0.01*3;
////assign chan_coeffs[19] = 0.01*3;

`else
output  rxp_out;

assign rxp_out = rx_in;

`endif


endmodule


//systemVerilog HDL for "wmu_lpddr4x_lib", "lpddr4x_nmos_switch" "systemVerilog"

`timescale 1ps/1fs
module wphy_sa_4g_2ph_pdly_no_esd_wphy_nmos_switch ( inn, inp, vss, ena, out);

`ifdef WPIN_EN
  input var integer inp;
  input var integer inn;
`else
  input inp;
  input inn;
`endif
  input ena;
  inout vss;
  output var integer out;

`ifdef WPIN_EN
`elsif WPIN_UART_EN
Wpin_uart_rx Winn(inn);
`endif


  wire pwr_ok;
  assign pwr_ok= ~vss;

`ifdef WCHANNEL_EN  var real `else logic `endif inp_channel;

wphy_sa_4g_2ph_pdly_no_esd_wphy_real_channel_model #(
     //parameters
     .COEFF_FILE         ( "channel_coeffs_10ps.txt"),
     .TIMESTEP_PS        ( 7        ),
     .NUM_OF_COEFFS      ( 20        ),
     .DELAY              ( 0        ),         // in ps
     .AMP_RATIO          ( 1        )         // 0<=value<=1,
   ) CH_00 (
     .rx_in(inp),
     .rxp_out(inp_channel));

 
`ifdef WPIN_EN 
  always @(*) begin
  	if (ena) begin
		if (inp === 32'bz) out = inn;
		else out = 32'bx;
	end
	else out = inp;
  
  end
  always @(*) begin
	if (~pwr_ok) out = 32'bx;
  end
`else
  always @(*) begin
  	if (ena) begin
`ifdef WPIN_UART_EN
		if (inp === 1'bz) out = Winn.value;
`else
		if (inp === 1'bz) out = inn*500;
`endif
		else out = 32'bx;
	end
	else out = inp_channel*1000;
  
  end
  always @(*) begin
	if (~pwr_ok) out = 32'bx;
  end
`endif


endmodule
`endif //SYNTHESIS
