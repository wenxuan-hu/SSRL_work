module crossbar_2ports_wrapper(
    input clk,rst,
    input [7:0] crb_READ_LATENCY_cfg,
    input [7:0] crb_WRITE_LATENCY_cfg,
    native_interface native_if_0,native_if_1,
    litedram_interface litedram_if
);
    crossbar_2ports u_crossbar_2ports (
    .interface_bank0_valid          (litedram_if.litedram_cmd_if_0.interface_bank_valid),
    .interface_bank0_ready          (litedram_if.litedram_cmd_if_0.interface_bank_ready),
    .interface_bank0_mw             (litedram_if.litedram_cmd_if_0.interface_bank_mw),
    .interface_bank0_we             (litedram_if.litedram_cmd_if_0.interface_bank_we),
    .interface_bank0_addr           (litedram_if.litedram_cmd_if_0.interface_bank_addr),
    .interface_bank0_lock           (litedram_if.litedram_cmd_if_0.interface_bank_lock),
    .interface_bank0_wdata_ready    (litedram_if.litedram_cmd_if_0.interface_bank_wdata_ready),
    .interface_bank0_rdata_valid    (litedram_if.litedram_cmd_if_0.interface_bank_rdata_valid),
    .interface_bank1_valid          (litedram_if.litedram_cmd_if_1.interface_bank_valid),
    .interface_bank1_ready          (litedram_if.litedram_cmd_if_1.interface_bank_ready),
    .interface_bank1_mw             (litedram_if.litedram_cmd_if_1.interface_bank_mw),
    .interface_bank1_we             (litedram_if.litedram_cmd_if_1.interface_bank_we),
    .interface_bank1_addr           (litedram_if.litedram_cmd_if_1.interface_bank_addr),
    .interface_bank1_lock           (litedram_if.litedram_cmd_if_1.interface_bank_lock),
    .interface_bank1_wdata_ready    (litedram_if.litedram_cmd_if_1.interface_bank_wdata_ready),
    .interface_bank1_rdata_valid    (litedram_if.litedram_cmd_if_1.interface_bank_rdata_valid),
    .interface_bank2_valid          (litedram_if.litedram_cmd_if_2.interface_bank_valid),
    .interface_bank2_ready          (litedram_if.litedram_cmd_if_2.interface_bank_ready),
    .interface_bank2_mw             (litedram_if.litedram_cmd_if_2.interface_bank_mw),
    .interface_bank2_we             (litedram_if.litedram_cmd_if_2.interface_bank_we),
    .interface_bank2_addr           (litedram_if.litedram_cmd_if_2.interface_bank_addr),
    .interface_bank2_lock           (litedram_if.litedram_cmd_if_2.interface_bank_lock),
    .interface_bank2_wdata_ready    (litedram_if.litedram_cmd_if_2.interface_bank_wdata_ready),
    .interface_bank2_rdata_valid    (litedram_if.litedram_cmd_if_2.interface_bank_rdata_valid),
    .interface_bank3_valid          (litedram_if.litedram_cmd_if_3.interface_bank_valid),
    .interface_bank3_ready          (litedram_if.litedram_cmd_if_3.interface_bank_ready),
    .interface_bank3_mw             (litedram_if.litedram_cmd_if_3.interface_bank_mw),
    .interface_bank3_we             (litedram_if.litedram_cmd_if_3.interface_bank_we),
    .interface_bank3_addr           (litedram_if.litedram_cmd_if_3.interface_bank_addr),
    .interface_bank3_lock           (litedram_if.litedram_cmd_if_3.interface_bank_lock),
    .interface_bank3_wdata_ready    (litedram_if.litedram_cmd_if_3.interface_bank_wdata_ready),
    .interface_bank3_rdata_valid    (litedram_if.litedram_cmd_if_3.interface_bank_rdata_valid),
    .interface_bank4_valid          (litedram_if.litedram_cmd_if_4.interface_bank_valid),
    .interface_bank4_ready          (litedram_if.litedram_cmd_if_4.interface_bank_ready),
    .interface_bank4_mw             (litedram_if.litedram_cmd_if_4.interface_bank_mw),
    .interface_bank4_we             (litedram_if.litedram_cmd_if_4.interface_bank_we),
    .interface_bank4_addr           (litedram_if.litedram_cmd_if_4.interface_bank_addr),
    .interface_bank4_lock           (litedram_if.litedram_cmd_if_4.interface_bank_lock),
    .interface_bank4_wdata_ready    (litedram_if.litedram_cmd_if_4.interface_bank_wdata_ready),
    .interface_bank4_rdata_valid    (litedram_if.litedram_cmd_if_4.interface_bank_rdata_valid),
    .interface_bank5_valid          (litedram_if.litedram_cmd_if_5.interface_bank_valid),
    .interface_bank5_ready          (litedram_if.litedram_cmd_if_5.interface_bank_ready),
    .interface_bank5_mw             (litedram_if.litedram_cmd_if_5.interface_bank_mw),
    .interface_bank5_we             (litedram_if.litedram_cmd_if_5.interface_bank_we),
    .interface_bank5_addr           (litedram_if.litedram_cmd_if_5.interface_bank_addr),
    .interface_bank5_lock           (litedram_if.litedram_cmd_if_5.interface_bank_lock),
    .interface_bank5_wdata_ready    (litedram_if.litedram_cmd_if_5.interface_bank_wdata_ready),
    .interface_bank5_rdata_valid    (litedram_if.litedram_cmd_if_5.interface_bank_rdata_valid),
    .interface_bank6_valid          (litedram_if.litedram_cmd_if_6.interface_bank_valid),
    .interface_bank6_ready          (litedram_if.litedram_cmd_if_6.interface_bank_ready),
    .interface_bank6_mw             (litedram_if.litedram_cmd_if_6.interface_bank_mw),
    .interface_bank6_we             (litedram_if.litedram_cmd_if_6.interface_bank_we),
    .interface_bank6_addr           (litedram_if.litedram_cmd_if_6.interface_bank_addr),
    .interface_bank6_lock           (litedram_if.litedram_cmd_if_6.interface_bank_lock),
    .interface_bank6_wdata_ready    (litedram_if.litedram_cmd_if_6.interface_bank_wdata_ready),
    .interface_bank6_rdata_valid    (litedram_if.litedram_cmd_if_6.interface_bank_rdata_valid),
    .interface_bank7_valid          (litedram_if.litedram_cmd_if_7.interface_bank_valid),
    .interface_bank7_ready          (litedram_if.litedram_cmd_if_7.interface_bank_ready),
    .interface_bank7_mw             (litedram_if.litedram_cmd_if_7.interface_bank_mw),
    .interface_bank7_we             (litedram_if.litedram_cmd_if_7.interface_bank_we),
    .interface_bank7_addr           (litedram_if.litedram_cmd_if_7.interface_bank_addr),
    .interface_bank7_lock           (litedram_if.litedram_cmd_if_7.interface_bank_lock),
    .interface_bank7_wdata_ready    (litedram_if.litedram_cmd_if_7.interface_bank_wdata_ready),
    .interface_bank7_rdata_valid    (litedram_if.litedram_cmd_if_7.interface_bank_rdata_valid),
    .interface_wdata                (litedram_if.litedram_data_if.interface_wdata),
    .interface_wdata_we             (litedram_if.litedram_data_if.interface_wdata_we),
    .interface_rdata                (litedram_if.litedram_data_if.interface_rdata),
    //csr
    .crb_READ_LATENCY_cfg           (crb_READ_LATENCY_cfg),
    .crb_WRITE_LATENCY_cfg          (crb_WRITE_LATENCY_cfg),
    //native0
    .cmd_valid                      (native_if_0.native_cmd_valid),
    .cmd_ready                      (native_if_0.native_cmd_ready),
    .cmd_first                      (native_if_0.native_cmd_first),
    .cmd_last                       (native_if_0.native_cmd_last),
    .cmd_payload_mw                 (native_if_0.native_cmd_payload_mw),
    .cmd_payload_we                 (native_if_0.native_cmd_payload_we),
    .cmd_payload_addr               (native_if_0.native_cmd_payload_addr),
    .wdata_valid                    (native_if_0.wdata_valid),
    .wdata_ready                    (native_if_0.wdata_ready),
    .wdata_first                    (native_if_0.wdata_first),
    .wdata_last                     (native_if_0.wdata_last),
    .wdata_payload_data             (native_if_0.wdata_payload_data),
    .wdata_payload_we               (native_if_0.wdata_payload_we),
    .rdata_valid                    (native_if_0.rdata_valid),
    .rdata_ready                    (native_if_0.rdata_ready),
    .rdata_first                    (native_if_0.rdata_first),
    .rdata_last                     (native_if_0.rdata_last),
    .rdata_payload_data             (native_if_0.rdata_payload_data),

    //native1
    .cmd_valid_1                    (native_if_1.native_cmd_valid),
    .cmd_ready_1                    (native_if_1.native_cmd_ready),
    .cmd_first_1                    (native_if_1.native_cmd_first),
    .cmd_last_1                     (native_if_1.native_cmd_last),
    .cmd_payload_mw_1               (native_if_1.native_cmd_payload_mw),
    .cmd_payload_we_1               (native_if_1.native_cmd_payload_we),
    .cmd_payload_addr_1             (native_if_1.native_cmd_payload_addr),
    .wdata_valid_1                  (native_if_1.wdata_valid),
    .wdata_ready_1                  (native_if_1.wdata_ready),
    .wdata_first_1                  (native_if_1.wdata_first),
    .wdata_last_1                   (native_if_1.wdata_last),
    .wdata_payload_data_1           (native_if_1.wdata_payload_data),
    .wdata_payload_we_1             (native_if_1.wdata_payload_we),
    .rdata_valid_1                  (native_if_1.rdata_valid),
    .rdata_ready_1                  (native_if_1.rdata_ready),
    .rdata_first_1                  (native_if_1.rdata_first),
    .rdata_last_1                   (native_if_1.rdata_last),
    .rdata_payload_data_1           (native_if_1.rdata_payload_data),
    .sys_clk                        (clk),
    .sys_rst                        (rst)
);
endmodule