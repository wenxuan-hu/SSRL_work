package bank_machine_test_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "tb_defs.svh"
    `include "bm_monitor.svh"

    `include "req_trans.svh"
    `include "req_cmd_sequence.svh"
    `include "req_sequencer.svh"
    `include "req_driver.svh"
    `include "req_monitor.svh"
    `include "req_agent.svh"

    `include "bm_responder.svh"
    `include "bank_machine_checker.svh"
    `include "bank_machine_virtual_sequencer.svh"
    `include "bank_machine_env.svh"
    `include "bank_machine_basic_test.svh"

endpackage